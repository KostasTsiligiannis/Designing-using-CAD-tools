module mlx (a, b, c, d, s, dp);
  input a, b, c, d;
  output [6:0] s;
  output         dp;
  wire[3:0] o;
  
  assign o = {a,b,c,d};
  assign s[6:0] = (o==4'b0000)? 7'b1110111: (o==4'b0001 )? 7'b0010010: (o==4'b0010) ? 7'b1011101 : (o==4'b0011)? 7'b1011011: (o==4'b0100) ? 7'b0111010 : (o==4'b0101) ? 7'b1101011 : (o==4'b0110) ? 7'b1101111 : (o==4'b0111) ? 7'b1011010 : (o==4'b1000) ? 7'b1111111 : (o==4'b1001) ? 7'b1111010 : (o==4'b1010) ? 7'b1111110 : (o==4'b1011) ? 7'b0101111 : (o==4'b1100) ? 7'b1100101 : (o==4'b1101) ? 7'b0011111 : (o==4'b1110) ? 7'b1101101 : (o==4'b1111) ? 7'b1101100 : 7'b0000000;
  assign dp = 1;
  
endmodule